module fifo (
	input clk,    // Clock
	
);

endmodule