module i2c_master
 (
 	input logic clk_in,
 	input logic reset_in,
 	input logic 
 	);
endmodule