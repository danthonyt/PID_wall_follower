module adc_lut_tb ();

endmodule