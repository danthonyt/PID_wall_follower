module top ();
// dc motor has time constant = 100ms
// pwm should be 100 Hz frequency
endmodule